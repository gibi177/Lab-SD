--Descrição: Implementação de um somador de palavras de 4 bits utilizando somadores completos

-- ****************************************** 
--  Circuito: Somador de palavras de 4 bits:
--  A Entrada 1
--  B Entrada 2
--  S Saida
-- ******************************************


-- Bibliotecas
library IEEE;
use ieee.std_logic_1164.ALL;

-- Entidade
entity Q1 is
    port (

    );
